`timescale 1ns/1ns
package agent_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;
    import dutb_param_pkg::*;
    import dutb_pkg::*;

    import dut_param_pkg::*;

    `include "dut_cin_driver.svh"
    // `include "dutb_pout_monitor.svh"
    // `include "dut_xds_in_driver.svh"
    // `include "dut_xds_out_driver.svh"
    // `include "dut_xds_in_frame_driver.svh"
    // `include "dut_xds_in_frame_monitor.svh"
    
endpackage
 