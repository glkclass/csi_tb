/******************************************************************************************************************************
    Project         :   CSI
    Creation Date   :   Dec 2021
    Interface       :   dut_if
    Description     :   
******************************************************************************************************************************/


// ****************************************************************************************************************************
interface dut_if(input 
                bit                     rst, hs_clk, csi_clk, 
                ci_if                   ci_vif, 
                fifo_if                 fifo_vif,
                d_phy_appi_if           d_phy_appi_vif,
                d_phy_adapter_line_if   d_phy_adapter_line_vif);
endinterface
// ****************************************************************************************************************************
