package scb_pkg;
    `include "uvm_macros.svh"
    // import uvm_pkg::*;
    import dutb_pkg::*;

endpackage
