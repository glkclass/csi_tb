`timescale 1ns/1ns
package test_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;

    import dutb_typedef_pkg::*;
    import dutb_pkg::*;
    
    import dut_param_pkg::*;
    import dut_if_proxy_pkg::*;
    import agent_pkg::*;
    import sequence_pkg::*;
    `include "dut_test.svh"
endpackage




