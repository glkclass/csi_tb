package scb_pkg;
    `include "uvm_macros.svh"
    // import uvm_pkg::*;
    import dut_scb_pkg::*;

endpackage
