`timescale 1ns/1ns
package test_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;
    import dut_test_pkg::*;

    import typedef_pkg::*;
    import dut_tb_param_pkg::*;
    import dut_handler_pkg::*;
    import dut_env_pkg::*;
    import agent_pkg::*;
    import dut_scb_pkg::*;
    import sequence_pkg::*;
    `include "dut_test.svh"


endpackage




