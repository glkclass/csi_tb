package dut_if_proxy_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;

    import dutb_pkg::*;
    `include "dut_if_proxy.svh"
endpackage


 
 
